BZh91AY&SYu�� _�Py�_�g߰?���P^t�F���Jx�L�F�� 1��&�R����2h2h�d 24ɦ� �LL%4(iM�&�P   ��&d`bba0�!�&�	M5d�@L!�=�~���h��	�$�I��f�
L��0�&�}F��ƀm�Si/	�����Z�m��F������8}�S�Ce�Fc��V�-$�i�-��ڠ�,h� JS��Z��|���'�r�2&=ҳj]1����@�L d6Zmƾ`�0�u3$�R$�s�S�C��<[9J*�-�w���C`B*	!!ƶ����]qz�h���2�H�'Ft�T��CAђ]�H�d��Ӵ��5����e*W��:ʾ�]	��'�� b���y�0��.
@�#�E��*�e<�Fcw���QP>kb8ٸ��i���3�mר�>�*���rJ=�F�"�!(�&����W$)K=j|�F�"D��5E�}��0�0�C��NDd�����d��M����O�\��J�7� ����%�[�ȁ<ɮ:�xi��/ЪOU�%d�_�8ek^��(�-��\ֳ�.������bh��K�;��۸��h�x��-�1!e�j%x� 6�<u�#ߐ�H&��!&ϖB�Q�h+v��D&װ����
�<-=�!�ar��S�w+�b ��[�p3A�s�kg4,�w�fԃzlZ���zk+X�Ic
��������쐈*ct��-�0�E@	(\��_���D�!Z$�e�#����\�i��Y��@j��Ɨ̽V�1y�6#rE����rE8P�u��